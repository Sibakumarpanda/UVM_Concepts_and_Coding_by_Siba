Example9: for set_type_override_by_type with parameterized classes
Note: For parameterized classes, an overriding class should have the same parameter values.
