Factory Overriding:
Based on the requirement, the behavior of the testbench can be changed by substituting one class with another when it is constructed. 
It is the process that allows an object of one type to be overridden with an object of its derived type without changing the testbench structure.   
This facility of the uvm factory allows users to override the class without editing or recompiling the code.
