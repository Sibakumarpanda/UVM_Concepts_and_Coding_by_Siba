Sequence-Driver-Sequencer communication in UVM :
-We discussed sequece_item, sequence, sequencer, and driver independently. 
-In this section, we will discuss how they talk with each other and provide sequence items from sequence to driver via the sequencer. 
-Before you start reading this section, make sure you are aware of all methods used in sequencer and driver. (Refer: UVM Sequencer and UVM Driver).
