Example1: Using get_next_item and item_done methods in the driver (Without RSP packet )
