uvm_resource_db in UVM:

-The uvm_resource_db is a type-parameterized class that is a convenience layer on the top of a resource database. 
-This convenience layer provides simplified access to the low-level database and it adds no new functionality. 
-Hence, uvm_resource_db is not derived from the uvm_resource class. 
-The below code snippet for the uvm_resource_db class is taken from the uvm source code.
