UVM Heartbeat example: Fail case
  
