UVM Heartbeat Example1: Success case
