Example10: for set_type_override_by_type with parameterized classes (with Different parameter)
Note: For parameterized classes, an overriding class should have the same parameter values.
      If an overriding class has different parameter values, factory overriding will fail.
