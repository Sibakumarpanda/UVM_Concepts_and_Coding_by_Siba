UVM Printer Understanding:
-The uvm_printer class provides flexibility to print uvm_objects in different formats. 
-We have discussed the print() method using `uvm_field_* macro or write do_print() method if utils_begin/ end macros are not used.
-The UVM printer provides four built-in printers.
  1.uvm_printer
  2.uvm_table_printer
  3.uvm_tree_printer
  4.uvm_line_printer
