UVM Heartbeat Concept Understanding:
