Example2: Using get_next_item and item_done methods in the driver (RSP packet)
