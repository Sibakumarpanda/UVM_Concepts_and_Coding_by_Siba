Example4: set_auto_reset method example
