//Example2: Example of Two agent uses with using Virtual Sequence and without Virtual Sequencer concept
