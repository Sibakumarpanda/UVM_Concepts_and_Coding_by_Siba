Example2: reset, get_threshold, and get_num_waiters methods example
