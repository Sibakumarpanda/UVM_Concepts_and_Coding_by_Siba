Example3: Using get and put methods in driver
