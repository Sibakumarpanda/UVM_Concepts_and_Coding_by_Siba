UVM Object:

The uvm_object class is the base class for all uvm hierarchical classes such as uvm_report_object, uvm_component, uvm_transaction, uvm_sequence_item, uvm_sequence etc. 
It serves an important role to define a set of methods such as create, copy, print, clone, compare, record, etc.

UVM Utility Macros and field macros:
