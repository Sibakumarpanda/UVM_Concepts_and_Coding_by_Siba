Example3: cancel method example
