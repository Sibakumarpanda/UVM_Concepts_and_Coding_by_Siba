UVM Heartbeat example:(With multiple components)
