Arbitration in Sequencer:
-The uvm_sequencer has a built-in mechanism to arbitrate within concurrently running sequences over the sequencer. 
-Based on the arbitration algorithm, the sequencer sends sequence_item to the driver for the granted sequence.
