Example9: for set_type_override_by_type with parameterized classes (same parameter)
Note: For parameterized classes, an overriding class should have the same parameter values, else it will fail.
